module x; a (x,y,.z(q); endmodule
     module y;
	     input a;
	     a
	        (.aa(aa),
		 .bb(bb))
	     ;
`define FOO 11
`ifdef FOO
	     b
	     (cin)
	     ;
`endif
	     endmodule
