module x;
a a (x, // commant
    y  /*com
	ment*/,
   .z(q);
endmodule
